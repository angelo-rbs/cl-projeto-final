library IEEE;
use IEEE.std_logic_1164.all;


ENTITY hex_to_seg_decoder IS
PORT (
	x0: IN STD_LOGIC;
	x1: IN STD_LOGIC;
	x2: IN STD_LOGIC;
	x3: IN STD_LOGIC;

	a: IN STD_LOGIC;
	b: IN STD_LOGIC;
	c: IN STD_LOGIC;
	d: IN STD_LOGIC;
	e: IN STD_LOGIC;
	f: IN STD_LOGIC;
	g: IN STD_LOGIC

     );
END hex_to_seg_decoder;

ARCHITECTURE impl OF hex_to_seg_decoder IS
BEGIN

END impl;

