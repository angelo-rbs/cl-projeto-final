library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity projeto is
    generic (
        TAM_REG : integer := 16  -- Tamanho de cada registrador
    );
    port (
        clk         : in  std_logic;
        reset       : in  std_logic;
        entrada     : in std_logic_vector(TAM_REG-1 downto 0);

        display        : out  std_logic_vector(0 to 27); -- valor atual
        display_estado : out std_logic_vector(0 to 6); -- estado atual

        ler_a       : in std_logic;
        ler_b       : in std_logic;
        calcular    : in std_logic
    );
end projeto;

architecture behaviour of projeto is

    component hex_to_seg is 
        port (
            entry: IN std_logic_vector(3 downto 0);
            segs: OUT std_logic_vector(0 to 6)
        );
    end component;

    component banco is 
        generic (
            NUM : integer := 8;  -- Número de registradores
            TAM_REG : integer := 16  -- Tamanho de cada registrador
        );
        port (
            clk         : in  std_logic;
            reset       : in  std_logic;
            entrada     : in std_logic_vector(TAM_REG-1 downto 0);
            saida       : out std_logic_vector(TAM_REG-1 downto 0);
            set_reg     : in  std_logic;
            set_val     : in  std_logic;
            get_val     : in  std_logic
        );
    end component;

    -- Estados gerais
    signal visor       : std_logic_vector(15 downto 0) := (others => '0');
    signal codigo_estado_em_binario : std_logic_vector(3 downto 0) := "1010";
    signal saida_banco : std_logic_vector(15 downto 0);

    -- Estados da divisão
    signal quoc : signed(15 downto 0) := (others => '0');
    signal dividendo : signed(15 downto 0) := (others => '0');
    signal divisor : signed(15 downto 0) := (others => '0');
    signal temp : signed(15 downto 0) := (others => '0');  -- Auxiliar para o loop de divisão
    
    -- Estados de entrada
    signal entrada_var   : std_logic_vector(TAM_REG-1 downto 0) := (others => '0');
    signal entrada_banco : std_logic_vector(TAM_REG-1 downto 0) := (others => '0');
    
    -- Estados de saída
    signal set_reg_control : std_logic := '0';
    signal set_val_control : std_logic := '0';
    signal get_val_control : std_logic := '1';

    -- Estado de controle para a divisão
    type state_type is (IDLE, READ_A, READ_B, DIVIDE, DONE);
    signal state, next_state : state_type := IDLE;

begin

    -- Instâncias dos componentes
    seg_a : hex_to_seg port map(
        entry => entrada_var(3 downto 0),
        segs => display(0 to 6)
    );
    seg_b : hex_to_seg port map(
        entry => entrada_var(7 downto 4),
        segs => display(7 to 13)
    );
    seg_c : hex_to_seg port map(
        entry => entrada_var(11 downto 8),
        segs => display(14 to 20)
    );
    seg_d : hex_to_seg port map(
        entry => entrada_var(15 downto 12),
        segs => display(21 to 27)
    );
    seg_estado : hex_to_seg port map(
        entry => codigo_estado_em_binario,
        segs => display_estado
    );
    
    banco_impl: banco 
    port map(
        clk => clk,
        reset => reset,
        entrada => entrada_banco,
        saida => saida_banco,
        set_reg => set_reg_control,
        set_val => set_val_control,
        get_val => get_val_control
    );

    -- Processo de controle de estado
    process(clk, reset)
    begin
        if reset = '0' then
            state <= IDLE;
            codigo_estado_em_binario <= "1010";
            entrada_banco <= (others => '0');
            set_reg_control <= '1';
            set_val_control <= '1';
            get_val_control <= '0';
            quoc <= (others => '0');
            dividendo <= (others => '0');
            divisor <= (others => '0');
            entrada_var <= (others => '0');
        elsif rising_edge(clk) then
            state <= next_state;
            
            case state is
                when IDLE =>
                    if ler_a = '0' then
                        next_state <= READ_A;
                    elsif ler_b = '0' then
                        next_state <= READ_B;
                    elsif calcular = '0' then
                        next_state <= DIVIDE;
                    else
                        next_state <= IDLE;
                    end if;
                    
                when READ_A =>
                    codigo_estado_em_binario <= "1010";
                    entrada_banco <= "0000000000000000";
                    set_reg_control <= '0';
                    set_val_control <= '1';
                    get_val_control <= '1';
                    next_state <= IDLE;
                    if get_val_control = '1' then
                        dividendo <= signed(saida_banco);
                    end if;
                    
                when READ_B =>
                    codigo_estado_em_binario <= "1011";
                    entrada_banco <= "0000000000000001";
                    set_reg_control <= '1';
                    set_val_control <= '0';
                    get_val_control <= '0';
                    next_state <= IDLE;
                    if get_val_control = '1' then
                        divisor <= signed(saida_banco);
                    end if;
                    
                when DIVIDE =>
                    codigo_estado_em_binario <= "1100";
                    quoc <= (others => '0');
                    temp <= dividendo;
                    
                    -- Divisão usando abordagem de subtração repetida
                    if temp >= divisor then
                        temp <= temp - divisor;
                        quoc <= quoc + 1;
                    else
                        next_state <= DONE;
                    end if;
                    
                when DONE =>
                    entrada_var <= std_logic_vector(quoc);
                    next_state <= IDLE;
                    
                when others =>
                    next_state <= IDLE;
            end case;
        end if;
    end process;
end behaviour;
